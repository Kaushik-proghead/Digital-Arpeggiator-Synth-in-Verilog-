// dds.v
`timescale 1ns/1ps
module dds #(
    parameter PHASE_WIDTH = 32,
    parameter OUT_WIDTH = 16,
    parameter LUT_ADDR_BITS = 8
)(
    input clk,
    input rst,
    input [PHASE_WIDTH-1:0] delta,   // step size; delta==0 => REST (silence)
    input [1:0] wave_sel,            // 00=sine, 01=square, 10=triangle, 11=saw
    output reg signed [OUT_WIDTH-1:0] out_sample
);

    reg [PHASE_WIDTH-1:0] phase;

    localparam LUT_SIZE = (1 << LUT_ADDR_BITS);
    reg signed [OUT_WIDTH-1:0] sine_rom [0:LUT_SIZE-1];

    initial begin
        // file generated by generate_sine_mem.py
        $readmemh("sine256.mem", sine_rom);
    end

    wire [LUT_ADDR_BITS-1:0] addr = phase[PHASE_WIDTH-1 -: LUT_ADDR_BITS];

    // rough saw and triangle derived from phase MSBs (simple)
    wire [OUT_WIDTH-1:0] top_bits_for_shape = phase[PHASE_WIDTH-1 -: OUT_WIDTH];
    wire signed [OUT_WIDTH-1:0] saw_val = {top_bits_for_shape};
    // triangle: map top N bits into triangular shape
    reg signed [OUT_WIDTH-1:0] tri_val;
    always @(*) begin
        // reflect the top 9 bits to make triangle-like shape (approx)
        if (phase[PHASE_WIDTH-1 -: (LUT_ADDR_BITS+1)] < (1 << LUT_ADDR_BITS))
            tri_val = top_bits_for_shape;
        else
            tri_val = -top_bits_for_shape;
    end

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            phase <= 0;
            out_sample <= 0;
        end else begin
            if (delta == 0) begin
                // REST: produce silence, don't advance phase
                out_sample <= 0;
            end else begin
                phase <= phase + delta;
                case (wave_sel)
                    2'b00: out_sample <= sine_rom[addr];
                    2'b01: out_sample <= (phase[PHASE_WIDTH-1] ? -16'sh7FFF : 16'sh7FFF);
                    2'b10: out_sample <= tri_val;
                    2'b11: out_sample <= saw_val;
                    default: out_sample <= sine_rom[addr];
                endcase
            end
        end
    end
endmodule
